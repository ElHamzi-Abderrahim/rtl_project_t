`ifndef OTHER_PKGS_SV
`define OTHER_PKGS_SV

	// `include "macros.svh"
	// `include "some_other_pkgs_fname.svh"

    package other_pkgs;
        // import uvm_pkg::* ;
        // import some_other_pkgs::* ;
        
        // `include "other_includes.sv"
		
    endpackage

`endif // `ifndef OTHER_PKGS_SV
