`include "dummy_module.v"