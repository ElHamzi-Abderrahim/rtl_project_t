`ifndef TB_DEFINES_SV
`define TB_DEFINES_SV

    `ifndef PARAM_VALUE
        `define PARAM_VALUE 7
    `endif


`endif
